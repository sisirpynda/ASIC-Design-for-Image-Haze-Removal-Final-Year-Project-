module lut(number,inverse);
 input [7:0] number;
 output reg [11:0] inverse;

always @(number)
begin
case(number)

8'b00000001 : inverse = 12'b111111111111;
8'b00000010 : inverse = 12'b100000000000;
8'b00000011 : inverse = 12'b010101010101;
8'b00000100 : inverse = 12'b010000000000;
8'b00000101 : inverse = 12'b001100110011;
8'b00000110 : inverse = 12'b001010101010;
8'b00000111 : inverse = 12'b001001001001;
8'b00001000 : inverse = 12'b001000000000;
8'b00001001 : inverse = 12'b000111000111;
8'b00001010 : inverse = 12'b000110011001;
8'b00001011 : inverse = 12'b000101110100;
8'b00001100 : inverse = 12'b000101010101;
8'b00001101 : inverse = 12'b000100111011;
8'b00001110 : inverse = 12'b000100100100;
8'b00001111 : inverse = 12'b000100010001;
8'b00010000 : inverse = 12'b000100000000;
8'b00010001 : inverse = 12'b000011110000;
8'b00010010 : inverse = 12'b000011100011;
8'b00010011 : inverse = 12'b000011010111;
8'b00010100 : inverse = 12'b000011001100;
8'b00010101 : inverse = 12'b000011000011;
8'b00010110 : inverse = 12'b000010111010;
8'b00010111 : inverse = 12'b000010110010;
8'b00011000 : inverse = 12'b000010101010;
8'b00011001 : inverse = 12'b000010100011;
8'b00011010 : inverse = 12'b000010011101;
8'b00011011 : inverse = 12'b000010010111;
8'b00011100 : inverse = 12'b000010010010;
8'b00011101 : inverse = 12'b000010001101;
8'b00011110 : inverse = 12'b000010001000;
8'b00011111 : inverse = 12'b000010000100;
8'b00100000 : inverse = 12'b000010000000;
8'b00100001 : inverse = 12'b000001111100;
8'b00100010 : inverse = 12'b000001111000;
8'b00100011 : inverse = 12'b000001110101;
8'b00100100 : inverse = 12'b000001110001;
8'b00100101 : inverse = 12'b000001101110;
8'b00100110 : inverse = 12'b000001101011;
8'b00100111 : inverse = 12'b000001101001;
8'b00101000 : inverse = 12'b000001100110;
8'b00101001 : inverse = 12'b000001100011;
8'b00101010 : inverse = 12'b000001100001;
8'b00101011 : inverse = 12'b000001011111;
8'b00101100 : inverse = 12'b000001011101;
8'b00101101 : inverse = 12'b000001011011;
8'b00101110 : inverse = 12'b000001011001;
8'b00101111 : inverse = 12'b000001010111;
8'b00110000 : inverse = 12'b000001010101;
8'b00110001 : inverse = 12'b000001010011;
8'b00110010 : inverse = 12'b000001010001;
8'b00110011 : inverse = 12'b000001010000;
8'b00110100 : inverse = 12'b000001001110;
8'b00110101 : inverse = 12'b000001001101;
8'b00110110 : inverse = 12'b000001001011;
8'b00110111 : inverse = 12'b000001001010;
8'b00111000 : inverse = 12'b000001001001;
8'b00111001 : inverse = 12'b000001000111;
8'b00111010 : inverse = 12'b000001000110;
8'b00111011 : inverse = 12'b000001000101;
8'b00111100 : inverse = 12'b000001000100;
8'b00111101 : inverse = 12'b000001000011;
8'b00111110 : inverse = 12'b000001000010;
8'b00111111 : inverse = 12'b000001000001;
8'b01000000 : inverse = 12'b000001000000;
8'b01000001 : inverse = 12'b000000111111;
8'b01000010 : inverse = 12'b000000111110;
8'b01000011 : inverse = 12'b000000111101;
8'b01000100 : inverse = 12'b000000111100;
8'b01000101 : inverse = 12'b000000111011;
8'b01000110 : inverse = 12'b000000111010;
8'b01000111 : inverse = 12'b000000111001;
8'b01001000 : inverse = 12'b000000111000;
8'b01001001 : inverse = 12'b000000111000;
8'b01001010 : inverse = 12'b000000110111;
8'b01001011 : inverse = 12'b000000110110;
8'b01001100 : inverse = 12'b000000110101;
8'b01001101 : inverse = 12'b000000110101;
8'b01001110 : inverse = 12'b000000110100;
8'b01001111 : inverse = 12'b000000110011;
8'b01010000 : inverse = 12'b000000110011;
8'b01010001 : inverse = 12'b000000110010;
8'b01010010 : inverse = 12'b000000110001;
8'b01010011 : inverse = 12'b000000110001;
8'b01010100 : inverse = 12'b000000110000;
8'b01010101 : inverse = 12'b000000110000;
8'b01010110 : inverse = 12'b000000101111;
8'b01010111 : inverse = 12'b000000101111;
8'b01011000 : inverse = 12'b000000101110;
8'b01011001 : inverse = 12'b000000101110;
8'b01011010 : inverse = 12'b000000101101;
8'b01011011 : inverse = 12'b000000101101;
8'b01011100 : inverse = 12'b000000101100;
8'b01011101 : inverse = 12'b000000101100;
8'b01011110 : inverse = 12'b000000101011;
8'b01011111 : inverse = 12'b000000101011;
8'b01100000 : inverse = 12'b000000101010;
8'b01100001 : inverse = 12'b000000101010;
8'b01100010 : inverse = 12'b000000101001;
8'b01100011 : inverse = 12'b000000101001;
8'b01100100 : inverse = 12'b000000101000;
8'b01100101 : inverse = 12'b000000101000;
8'b01100110 : inverse = 12'b000000101000;
8'b01100111 : inverse = 12'b000000100111;
8'b01101000 : inverse = 12'b000000100111;
8'b01101001 : inverse = 12'b000000100111;
8'b01101010 : inverse = 12'b000000100110;
8'b01101011 : inverse = 12'b000000100110;
8'b01101100 : inverse = 12'b000000100101;
8'b01101101 : inverse = 12'b000000100101;
8'b01101110 : inverse = 12'b000000100101;
8'b01101111 : inverse = 12'b000000100100;
8'b01110000 : inverse = 12'b000000100100;
8'b01110001 : inverse = 12'b000000100100;
8'b01110010 : inverse = 12'b000000100011;
8'b01110011 : inverse = 12'b000000100011;
8'b01110100 : inverse = 12'b000000100011;
8'b01110101 : inverse = 12'b000000100011;
8'b01110110 : inverse = 12'b000000100010;
8'b01110111 : inverse = 12'b000000100010;
8'b01111000 : inverse = 12'b000000100010;
8'b01111001 : inverse = 12'b000000100001;
8'b01111010 : inverse = 12'b000000100001;
8'b01111011 : inverse = 12'b000000100001;
8'b01111100 : inverse = 12'b000000100001;
8'b01111101 : inverse = 12'b000000100000;
8'b01111110 : inverse = 12'b000000100000;
8'b01111111 : inverse = 12'b000000100000;
8'b10000000 : inverse = 12'b000000100000;
8'b10000001 : inverse = 12'b000000011111;
8'b10000010 : inverse = 12'b000000011111;
8'b10000011 : inverse = 12'b000000011111;
8'b10000100 : inverse = 12'b000000011111;
8'b10000101 : inverse = 12'b000000011110;
8'b10000110 : inverse = 12'b000000011110;
8'b10000111 : inverse = 12'b000000011110;
8'b10001000 : inverse = 12'b000000011110;
8'b10001001 : inverse = 12'b000000011101;
8'b10001010 : inverse = 12'b000000011101;
8'b10001011 : inverse = 12'b000000011101;
8'b10001100 : inverse = 12'b000000011101;
8'b10001101 : inverse = 12'b000000011101;
8'b10001110 : inverse = 12'b000000011100;
8'b10001111 : inverse = 12'b000000011100;
8'b10010000 : inverse = 12'b000000011100;
8'b10010001 : inverse = 12'b000000011100;
8'b10010010 : inverse = 12'b000000011100;
8'b10010011 : inverse = 12'b000000011011;
8'b10010100 : inverse = 12'b000000011011;
8'b10010101 : inverse = 12'b000000011011;
8'b10010110 : inverse = 12'b000000011011;
8'b10010111 : inverse = 12'b000000011011;
8'b10011000 : inverse = 12'b000000011010;
8'b10011001 : inverse = 12'b000000011010;
8'b10011010 : inverse = 12'b000000011010;
8'b10011011 : inverse = 12'b000000011010;
8'b10011100 : inverse = 12'b000000011010;
8'b10011101 : inverse = 12'b000000011010;
8'b10011110 : inverse = 12'b000000011001;
8'b10011111 : inverse = 12'b000000011001;
8'b10100000 : inverse = 12'b000000011001;
8'b10100001 : inverse = 12'b000000011001;
8'b10100010 : inverse = 12'b000000011001;
8'b10100011 : inverse = 12'b000000011001;
8'b10100100 : inverse = 12'b000000011000;
8'b10100101 : inverse = 12'b000000011000;
8'b10100110 : inverse = 12'b000000011000;
8'b10100111 : inverse = 12'b000000011000;
8'b10101000 : inverse = 12'b000000011000;
8'b10101001 : inverse = 12'b000000011000;
8'b10101010 : inverse = 12'b000000011000;
8'b10101011 : inverse = 12'b000000010111;
8'b10101100 : inverse = 12'b000000010111;
8'b10101101 : inverse = 12'b000000010111;
8'b10101110 : inverse = 12'b000000010111;
8'b10101111 : inverse = 12'b000000010111;
8'b10110000 : inverse = 12'b000000010111;
8'b10110001 : inverse = 12'b000000010111;
8'b10110010 : inverse = 12'b000000010111;
8'b10110011 : inverse = 12'b000000010110;
8'b10110100 : inverse = 12'b000000010110;
8'b10110101 : inverse = 12'b000000010110;
8'b10110110 : inverse = 12'b000000010110;
8'b10110111 : inverse = 12'b000000010110;
8'b10111000 : inverse = 12'b000000010110;
8'b10111001 : inverse = 12'b000000010110;
8'b10111010 : inverse = 12'b000000010110;
8'b10111011 : inverse = 12'b000000010101;
8'b10111100 : inverse = 12'b000000010101;
8'b10111101 : inverse = 12'b000000010101;
8'b10111110 : inverse = 12'b000000010101;
8'b10111111 : inverse = 12'b000000010101;
8'b11000000 : inverse = 12'b000000010101;
8'b11000001 : inverse = 12'b000000010101;
8'b11000010 : inverse = 12'b000000010101;
8'b11000011 : inverse = 12'b000000010101;
8'b11000100 : inverse = 12'b000000010100;
8'b11000101 : inverse = 12'b000000010100;
8'b11000110 : inverse = 12'b000000010100;
8'b11000111 : inverse = 12'b000000010100;
8'b11001000 : inverse = 12'b000000010100;
8'b11001001 : inverse = 12'b000000010100;
8'b11001010 : inverse = 12'b000000010100;
8'b11001011 : inverse = 12'b000000010100;
8'b11001100 : inverse = 12'b000000010100;
8'b11001101 : inverse = 12'b000000010011;
8'b11001110 : inverse = 12'b000000010011;
8'b11001111 : inverse = 12'b000000010011;
8'b11010000 : inverse = 12'b000000010011;
8'b11010001 : inverse = 12'b000000010011;
8'b11010010 : inverse = 12'b000000010011;
8'b11010011 : inverse = 12'b000000010011;
8'b11010100 : inverse = 12'b000000010011;
8'b11010101 : inverse = 12'b000000010011;
8'b11010110 : inverse = 12'b000000010011;
8'b11010111 : inverse = 12'b000000010011;
8'b11011000 : inverse = 12'b000000010010;
8'b11011001 : inverse = 12'b000000010010;
8'b11011010 : inverse = 12'b000000010010;
8'b11011011 : inverse = 12'b000000010010;
8'b11011100 : inverse = 12'b000000010010;
8'b11011101 : inverse = 12'b000000010010;
8'b11011110 : inverse = 12'b000000010010;
8'b11011111 : inverse = 12'b000000010010;
8'b11100000 : inverse = 12'b000000010010;
8'b11100001 : inverse = 12'b000000010010;
8'b11100010 : inverse = 12'b000000010010;
8'b11100011 : inverse = 12'b000000010010;
8'b11100100 : inverse = 12'b000000010001;
8'b11100101 : inverse = 12'b000000010001;
8'b11100110 : inverse = 12'b000000010001;
8'b11100111 : inverse = 12'b000000010001;
8'b11101000 : inverse = 12'b000000010001;
8'b11101001 : inverse = 12'b000000010001;
8'b11101010 : inverse = 12'b000000010001;
8'b11101011 : inverse = 12'b000000010001;
8'b11101100 : inverse = 12'b000000010001;
8'b11101101 : inverse = 12'b000000010001;
8'b11101110 : inverse = 12'b000000010001;
8'b11101111 : inverse = 12'b000000010001;
8'b11110000 : inverse = 12'b000000010001;
8'b11110001 : inverse = 12'b000000010000;
8'b11110010 : inverse = 12'b000000010000;
8'b11110011 : inverse = 12'b000000010000;
8'b11110100 : inverse = 12'b000000010000;
8'b11110101 : inverse = 12'b000000010000;
8'b11110110 : inverse = 12'b000000010000;
8'b11110111 : inverse = 12'b000000010000;
8'b11111000 : inverse = 12'b000000010000;
8'b11111001 : inverse = 12'b000000010000;
8'b11111010 : inverse = 12'b000000010000;
8'b11111011 : inverse = 12'b000000010000;
8'b11111100 : inverse = 12'b000000010000;
8'b11111101 : inverse = 12'b000000010000;
8'b11111110 : inverse = 12'b000000010000;
default : inverse = 12'b1111_1111_1111;
endcase 
end

endmodule

module test_lut;

reg [7:0] inn;
wire [11:0] outt;
wire [7:0]anss;

lut lt1(inn,outt);
assign anss = (outt*'d1000)>>12;

initial
begin
	inn = 'd250;
	#20
	inn = 'd200;
	#20
	inn = 'd100;
	#20
	inn = 'd50;
	#20
	inn = 'd10;
	#100 $finish;
end
endmodule  
